module RM_ctrl (
	input 						rst,
	input[`ByteSlctWidth-1:0]	byte_slct,
	input[`RegDataWidth-1:0]	raw_mem_data,

	output[`RegDataWidth-1:0]	data_to_reg
);
	//TODO
endmodule