module WM_ctrl (
	input 						rst,
	input[`RegDataWidth-1:0] 	raw_reg_data,
	input[`ByteSlctWidth-1:0]	byte_slct_MEM,

	output[`RegDataWidth-1:0]	data_to_mem
);
	// TODO
endmodule